-- Created on: 1993-01-18
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MaterialsDictionary from Materials 

	---Purpose: This class creates  a dictionary of materials.

inherits

    Transient
    
uses
    OStream           from  Standard,
    HAsciiString      from TCollection,
    MaterialsSequence from Materials,
    Material          from Materials

raises

    NoSuchObject from Standard

is

    Create returns mutable MaterialsDictionary from Materials;
    ---Level: Internal    
    ---Purpose: Returns a  MaterialsDictionary  object which  contains
    --          the sequence of all the   materials the user wants  to
    --          consider.
    
    Material(me ; amaterial : CString from Standard) returns Material from Materials    
    raises NoSuchObject from Standard   
    ---Level: Internal   
    ---Purpose: Retrieves from the dictionary the object material with
    --          <amaterial> as name.  If <amaterial> does not exist in
    --          the dictionary an exeption is raised.
    is static;
    
    ExistMaterial(me ; aName : CString from Standard) returns Boolean from Standard;
    ---Purpose: True if the materialofname aName exists ...
    
    NumberOfMaterials(me) returns Integer from Standard  
    ---Level: Internal 
    ---Purpose: Returns  the number of  materials previously stored in
    --          the dictionary.
    is static;
    
    Material(me ; anindex : Integer from Standard) returns Material from Materials
    ---Level: Internal
    ---Purpose: This method used  with  the  previous one, allow   the
    --          exploration  of   all  the  dictionary.  It  returns a
    --          Material instance.
    is static;
    
    UpToDate(me) returns Boolean from Standard
    ---Level: Internal
    ---Purpose: Returns true if there has been no  modification of the
    --          file Materials.dat  since the   creation of the dictionary
    --          object, false otherwise.  
    is static;
    
    Dump(me ; astream : in out OStream from Standard )
    ---Level: Internal
    ---Purpose: Useful for debugging.
    is static;
    
fields

    thefilename          : HAsciiString from TCollection;
    thetime              : Time from Standard;
    thematerialssequence : MaterialsSequence from Materials;

end MaterialsDictionary;
