-- Created on: 1992-02-18
-- Created by: Christophe MARION
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PolyAlgo from HLRBRep inherits TShared from MMgt

	---Purpose: to remove Hidden lines on Shapes with Triangulations.
      -- A framework to compute the shape as seen in
    	-- a projection plane. This is done by calculating
    	-- the visible and the hidden parts of the shape.
    	-- HLRBRep_PolyAlgo works with three types of entity:
    	-- -   shapes to be visualized (these shapes must
    	--   have already been triangulated.)
    	-- -   edges in these shapes (these edges are
    	--   defined as polygonal lines on the
    	--   triangulation of the shape, and are the basic
    	--   entities which will be visualized or hidden), and
    	-- -   triangles in these shapes which hide the edges.
    	--   HLRBRep_PolyAlgo is based on the principle
    	-- of comparing each edge of the shape to be
    	-- visualized with each of the triangles produced
    	-- by the triangulation of the shape, and
    	-- calculating the visible and the hidden parts of each edge.
    	-- For a given projection, HLRBRep_PolyAlgo
    	-- calculates a set of lines characteristic of the
    	-- object being represented. It is also used in
    	-- conjunction with the HLRBRep_PolyHLRToShape extraction
    	-- utilities, which reconstruct a new, simplified
    	-- shape from a selection of calculation results.
    	-- This new shape is made up of edges, which
    	-- represent the shape visualized in the projection.
    	-- HLRBRep_PolyAlgo works with a polyhedral
    	-- simplification of the shape whereas
    	-- HLRBRep_Algo takes the shape itself into
    	-- account. When you use HLRBRep_Algo, you
    	-- obtain an exact result, whereas, when you use
    	-- HLRBRep_PolyAlgo, you reduce computation
    	-- time but obtain polygonal segments.
    	-- An HLRBRep_PolyAlgo object provides a framework for:
    	-- -   defining the point of view
    	-- -   identifying the shape or shapes to be visualized
    	-- -   calculating the outlines
    	-- -   calculating the visible and hidden lines of the shape.
    	--   Warning
    	-- -   Superimposed lines are not eliminated by this algorithm.
    	-- -   There must be no unfinished objects inside the shape you wish to visualize.
    	-- -   Points are not treated.
    	-- -   Note that this is not the sort of algorithm
    	--   used in generating shading, which calculates
    	--   the visible and hidden parts of each face in a
    	--   shape to be visualized by comparing each
    	--   face in the shape with every other face in the same shape.

uses
    Address           from Standard,
    Boolean           from Standard,
    Integer           from Standard,
    Real              from Standard,
    Array1OfInteger   from TColStd,
    Array1OfTransient from TColStd,
    SequenceOfShape   from TopTools,
    IndexedMapOfShape from TopTools,
    MapOfShape        from TopTools,
    ListOfShape       from TopTools,
    Shape             from GeomAbs,
    Edge              from TopoDS,
    Shape             from TopoDS,
    Surface           from Geom,
    Curve2d           from BRepAdaptor,
    Curve             from BRepAdaptor,
    Surface           from BRepAdaptor,
    PolyInternalData  from HLRAlgo,
    ListOfBPoint      from HLRAlgo,
    TriangleData      from HLRAlgo,
    Projector         from HLRAlgo,
    EdgeStatus        from HLRAlgo,
    PolyAlgo          from HLRAlgo

raises
    OutOfRange   from Standard
    
is
    Create
    returns PolyAlgo from HLRBRep;
    	---Purpose: Constructs an empty framework for the
    	-- calculation of the visible and hidden lines of a shape in a projection.
    	-- Use the functions:
    	-- -   Projector to define the point of view
    	-- -   Load to select the shape or shapes to be  visualized
    	-- -   Update to compute the visible and hidden lines of the shape.
    	--   Warning
    	-- The shape or shapes to be visualized must have already been triangulated.
        
    Create(A : PolyAlgo from HLRBRep)
    returns PolyAlgo from HLRBRep;

    Create(S : Shape from TopoDS)
    returns PolyAlgo from HLRBRep;
    
    NbShapes(me) returns Integer from Standard
	---C++: inline
    is static;
    
    Shape(me : mutable; I : Integer from Standard)
    returns Shape from TopoDS
    raises OutOfRange from Standard
    	---C++: return &
    is static;
    
    Remove(me : mutable; I : Integer from Standard)
    raises OutOfRange from Standard
	---Purpose: remove the Shape of Index <I>.
    is static;

    Index(me; S : Shape from TopoDS) returns Integer from Standard
	---Purpose: return the index of the Shape <S> and  return 0 if
	--          the Shape <S> is not found.
    is static;

    Load(me : mutable; S : Shape from TopoDS)
	---Purpose: Loads the shape S into this framework.
    	-- Warning S must have already been triangulated.
   	---C++: inline
    	 is static;
    
    Algo(me) returns PolyAlgo from HLRAlgo
    is static;
    
    Projector(me) returns Projector from HLRAlgo
    	---Purpose: Sets the parameters of the view for this framework.
    	-- These parameters are defined by an HLRAlgo_Projector object,
    	-- which is returned by the Projector function on a Prs3d_Projector object.
        ---C++: return const &
	---C++: inline
    is static;
    
    Projector(me : mutable; P : Projector from HLRAlgo)
	---C++: inline
    is static;
    
    Angle(me) returns Real from Standard
	---C++: inline
    is static;
    
    Angle(me : mutable; Ang : Real from Standard)
	---C++: inline
    is static;
    
    TolAngular(me) returns Real from Standard
	---C++: inline
    is static;
    
    TolAngular(me : mutable; Tol : Real from Standard)
	---C++: inline
    is static;
    
    TolCoef(me) returns Real from Standard
	---C++: inline
    is static;
    
    TolCoef(me : mutable; Tol : Real from Standard)
	---C++: inline
    is static;
    
    Update(me : mutable)
	---Purpose: Launches calculation of outlines of the shape
    	-- visualized by this framework. Used after setting the point of view and
    	-- defining the shape or shapes to be visualized.
    is static;
    
    MakeShape(me) returns Shape from TopoDS
    is static private;

    InitShape(me      : mutable;
              Shape   :     Shape   from TopoDS;
	      IsoledF : out Boolean from Standard;
	      IsoledE : out Boolean from Standard)
    returns Integer from Standard
    is static private;

    StoreShell(me              : mutable;
               Shape           :     Shape             from TopoDS;
               iShell          : out Integer           from Standard;
               Shell           : out Array1OfTransient from TColStd;
	       IsoledF,IsoledE :     Boolean           from Standard; 
               ES              : out Array1OfInteger   from TColStd;
               PD,PID          : out Array1OfTransient from TColStd;
               ShapeMap1       : out MapOfShape        from TopTools;
               ShapeMap2       : out MapOfShape        from TopTools)
    is static private;
    
    Normal(me;
    	   iNode       :     Integer          from Standard;
           Nod1Indices :     Address          from Standard;
           Nod1RValues :     Address          from Standard;
	   TData       : out Address          from Standard;
	   PISeg       : out Address          from Standard;
	   PINod       : out Address          from Standard;
           orient      :     Boolean          from Standard) 
    returns Boolean from Standard
    is static private;
    
    AverageNormal(me; iNode       :     Integer from Standard;
                      Nod1Indices :     Address from Standard;
                      TData       : out Address from Standard;
                      PISeg       : out Address from Standard;
                      PINod       : out Address from Standard;
                      X,Y,Z       : out Real    from Standard)
    returns Boolean from Standard
    is static private;

    AddNormalOnTriangle(me; iTri  :     Integer from Standard;
                            iNode :     Integer from Standard;
                            jNode : out Integer from Standard;
                            TData : out Address from Standard;
                            PINod : out Address from Standard;
			    X,Y,Z : out Real    from Standard;
                            OK    : out Boolean from Standard)
    is static private;

    InitBiPointsWithConnexity
    	(me     : mutable;
         e      :     Integer           from Standard;
	 E      : out Edge              from TopoDS;
         List   : out ListOfBPoint      from HLRAlgo;
         PID    : out Array1OfTransient from TColStd;
	 LS     : out ListOfShape       from TopTools;
	 connex :     Boolean           from Standard)
    is static private;

    Interpolation(me;
                  List           : out ListOfBPoint     from HLRAlgo;
	          X1  ,Y1  ,Z1   : out Real             from Standard;
                  X2  ,Y2  ,Z2   : out Real             from Standard;
                  XTI1,YTI1,ZTI1 : out Real             from Standard;
                  XTI2,YTI2,ZTI2 : out Real             from Standard;
		  e              :     Integer          from Standard;
		  U1,U2          : out Real             from Standard;
                  Nod11Indices   : out Address          from Standard;
                  Nod11RValues   : out Address          from Standard;
                  Nod12Indices   : out Address          from Standard;
                  Nod12RValues   : out Address          from Standard;
		  i1p1,i1p2,i1   :     Integer          from Standard;
                  pid1           :     PolyInternalData from HLRAlgo;
                  TData1         : out Address          from Standard;
                  PISeg1         : out Address          from Standard;
		  PINod1         : out Address          from Standard)
    is static private;

    Interpolation(me;
                  List           : out ListOfBPoint     from HLRAlgo;
	          X1  ,Y1  ,Z1   : out Real             from Standard;
                  X2  ,Y2  ,Z2   : out Real             from Standard;
                  XTI1,YTI1,ZTI1 : out Real             from Standard;
                  XTI2,YTI2,ZTI2 : out Real             from Standard;
		  e              :     Integer          from Standard;
		  U1,U2          : out Real             from Standard;
		  rg             :     Shape            from GeomAbs;
                  Nod11Indices   : out Address          from Standard;
                  Nod11RValues   : out Address          from Standard;
                  Nod12Indices   : out Address          from Standard;
                  Nod12RValues   : out Address          from Standard;
		  i1p1,i1p2,i1   :     Integer          from Standard;
                  pid1           :     PolyInternalData from HLRAlgo;
                  TData1         : out Address          from Standard;
                  PISeg1         : out Address          from Standard;
		  PINod1         : out Address          from Standard;
                  Nod21Indices   : out Address          from Standard;
                  Nod21RValues   : out Address          from Standard;
                  Nod22Indices   : out Address          from Standard;
                  Nod22RValues   : out Address          from Standard;
		  i2p1,i2p2,i2   :     Integer          from Standard;
                  pid2           :     PolyInternalData from HLRAlgo;
                  TData2         : out Address          from Standard;
                  PISeg2         : out Address          from Standard;
		  PINod2         : out Address          from Standard)
    is static private;

    Interpolation(me;
		  U1,U2       :     Real    from Standard;
                  Nod1RValues :     Address from Standard;
                  Nod2RValues :     Address from Standard;
                  X3,Y3,Z3    : out Real    from Standard;
                  XT3,YT3,ZT3 : out Real    from Standard;
		  coef3,U3    : out Real    from Standard;
		  mP3P1       : out Boolean from Standard)
    returns Boolean from Standard
    is static private;

    MoveOrInsertPoint(me;
                      List           : out ListOfBPoint     from HLRAlgo;
                      X1  ,Y1  ,Z1   : out Real             from Standard;
                      X2  ,Y2  ,Z2   : out Real             from Standard;
                      XTI1,YTI1,ZTI1 : out Real             from Standard;
                      XTI2,YTI2,ZTI2 : out Real             from Standard;
		      e              :     Integer          from Standard;
		      U1,U2          : out Real             from Standard;
                      Nod11Indices   : out Address          from Standard;
                      Nod11RValues   : out Address          from Standard;
                      Nod12Indices   : out Address          from Standard;
                      Nod12RValues   : out Address          from Standard;
		      i1p1,i1p2,i1   :     Integer          from Standard;
                      pid1           :     PolyInternalData from HLRAlgo;
                      TData1         : out Address          from Standard;
                      PISeg1         : out Address          from Standard;
	              PINod1         : out Address          from Standard;
                      X3,Y3,Z3       :     Real             from Standard;
                      XT3,YT3,ZT3    :     Real             from Standard;
	              coef3          :     Real             from Standard;
	              U3             :     Real             from Standard;
                      insP3,mP3P1    :     Boolean          from Standard; 
		      flag           :     Integer          from Standard)
    is static private;

    MoveOrInsertPoint(me;
                      List           : out ListOfBPoint     from HLRAlgo;
                      X1  ,Y1  ,Z1   : out Real             from Standard;
                      X2  ,Y2  ,Z2   : out Real             from Standard;
                      XTI1,YTI1,ZTI1 : out Real             from Standard;
                      XTI2,YTI2,ZTI2 : out Real             from Standard;
		      e              :     Integer          from Standard;
		      U1,U2          : out Real             from Standard;
                      Nod11Indices   : out Address          from Standard;
                      Nod11RValues   : out Address          from Standard;
                      Nod12Indices   : out Address          from Standard;
                      Nod12RValues   : out Address          from Standard;
		      i1p1,i1p2,i1   :     Integer          from Standard;
                      pid1           :     PolyInternalData from HLRAlgo;
                      TData1         : out Address          from Standard;
                      PISeg1         : out Address          from Standard;
	              PINod1         : out Address          from Standard;
                      Nod21Indices   : out Address          from Standard;
                      Nod21RValues   : out Address          from Standard;
                      Nod22Indices   : out Address          from Standard;
                      Nod22RValues   : out Address          from Standard;
		      i2p1,i2p2,i2   :     Integer          from Standard;
                      pid2           :     PolyInternalData from HLRAlgo;
                      TData2         : out Address          from Standard;
                      PISeg2         : out Address          from Standard;
	              PINod2         : out Address          from Standard;
                      X3,Y3,Z3       :     Real             from Standard;
		      XT3,YT3,ZT3    :     Real             from Standard;
	              coef3          :     Real             from Standard;
	              U3             :     Real             from Standard;
                      insP3,mP3P1    :     Boolean          from Standard; 
		      flag           :     Integer          from Standard)
    is static private;

    MoveOrInsertPoint(me;
                      List           : out ListOfBPoint     from HLRAlgo;
                      X1  ,Y1  ,Z1   : out Real             from Standard;
                      X2  ,Y2  ,Z2   : out Real             from Standard;
                      XTI1,YTI1,ZTI1 : out Real             from Standard;
                      XTI2,YTI2,ZTI2 : out Real             from Standard;
		      e              :     Integer          from Standard;
		      U1,U2          : out Real             from Standard;
                      Nod11Indices   : out Address          from Standard;
                      Nod11RValues   : out Address          from Standard;
                      Nod12Indices   : out Address          from Standard;
                      Nod12RValues   : out Address          from Standard;
		      i1p1,i1p2,i1   :     Integer          from Standard;
                      pid1           :     PolyInternalData from HLRAlgo;
                      TData1         : out Address          from Standard;
                      PISeg1         : out Address          from Standard;
	              PINod1         : out Address          from Standard;
                      Nod21Indices   : out Address          from Standard;
                      Nod21RValues   : out Address          from Standard;
                      Nod22Indices   : out Address          from Standard;
                      Nod22RValues   : out Address          from Standard;
		      i2p1,i2p2,i2   :     Integer          from Standard;
                      pid2           :     PolyInternalData from HLRAlgo;
                      TData2         : out Address          from Standard;
                      PISeg2         : out Address          from Standard;
	              PINod2         : out Address          from Standard;
                      X3,Y3,Z3       :     Real             from Standard;
		      XT3,YT3,ZT3    :     Real             from Standard;
	              coef3          :     Real             from Standard;
	              U3             :     Real             from Standard;
                      insP3,mP3P1    :     Boolean          from Standard; 
                      X4,Y4,Z4       :     Real             from Standard;
		      XT4,YT4,ZT4    :     Real             from Standard;
	              coef4          :     Real             from Standard;
	              U4             :     Real             from Standard;
                      insP4,mP4P1    :     Boolean          from Standard; 
		      flag           :     Integer          from Standard)
    is static private;

    InsertOnOutLine(me  : mutable;
                    PID : out Array1OfTransient from TColStd)
    is static private;
    
    CheckFrBackTriangles(me   : mutable;
                         List : out ListOfBPoint      from HLRAlgo;
                         PID  : out Array1OfTransient from TColStd)
    is static private;
    
    FindEdgeOnTriangle(me;
		       Tri1Indices :     Address from Standard; 
	               ip1,ip2     :     Integer from Standard; 
                       jtrouv      : out Integer from Standard; 
                       isDirect    : out Boolean from Standard) 
    is static private;

    ChangeNode(me;
               ip1,ip2     :     Integer from Standard;
               Nod1Indices :     Address from Standard;
               Nod1RValues :     Address from Standard;
               Nod2Indices :     Address from Standard;
               Nod2RValues :     Address from Standard;
	       coef1       :     Real    from Standard;
               X3,Y3,Z3    :     Real    from Standard;
               first       :     Boolean from Standard;
               TData       : out Address from Standard;
               PISeg       : out Address from Standard;
               PINod       : out Address from Standard)
    is static private;
    
    UpdateAroundNode(me;
                     iNode       : Integer from Standard;
                     Nod1Indices : Address from Standard;
                     TData       : Address from Standard;
                     PISeg       : Address from Standard;
                     PINod       : Address from Standard)
    is static private;

    OrientTriangle(me ;iTri        : Integer from Standard;
                       Tri1Indices : Address from Standard;
                       Nod1Indices : Address from Standard;
                       Nod1RValues : Address from Standard;
                       Nod2Indices : Address from Standard;
                       Nod2RValues : Address from Standard;
                       Nod3Indices : Address from Standard;
                       Nod3RValues : Address from Standard)
    is static private;

    Triangles(me; ip1,ip2     :     Integer from Standard;
                  Nod1Indices :     Address from Standard;
                  PISeg       : out Address from Standard;
                  iTri1,iTri2 : out Integer from Standard)
    returns Boolean from Standard
    is static private;

    NewNode(me;
            Nod1RValues :     Address from Standard;
            Nod2RValues :     Address from Standard;
	    coef1       : out Real    from Standard;
            moveP1      : out Boolean from Standard)
    returns Boolean from Standard
    is static private;
    
    UVNode(me;
           Nod1RValues :     Address from Standard;
           Nod2RValues :     Address from Standard;
	   coef1       :     Real    from Standard;
           U3,V3       : out Real    from Standard)
    is static private;
    
    CheckDegeneratedSegment(me;
                            Nod1Indices : Address from Standard;
                            Nod1RValues : Address from Standard;
                            Nod2Indices : Address from Standard;
                            Nod2RValues : Address from Standard)
    is static private;

    UpdateOutLines(me   : mutable;
                   List : out ListOfBPoint      from HLRAlgo;
                   PID  : out Array1OfTransient from TColStd)
    is static private;
    
    UpdateEdgesBiPoints(me     : mutable;
                        List   : out ListOfBPoint      from HLRAlgo;
			PID    :     Array1OfTransient from TColStd;
                        closed :     Boolean           from Standard)
    is static private;
    
    UpdatePolyData(me     : mutable;
                   PD,PID : out Array1OfTransient from TColStd;
                   closed :     Boolean           from Standard)
    is static private;
    
    TMultiply(me;
              X,Y,Z : out Real from Standard;
              VecPartOnly : Boolean from Standard = Standard_False)
    is static private;
    
    TTMultiply(me;
               X,Y,Z : out Real from Standard;
              VecPartOnly : Boolean from Standard = Standard_False)
    is static private;
    
    TIMultiply(me;
               X,Y,Z : out Real from Standard;
               VecPartOnly : Boolean from Standard = Standard_False)
    is static private;
    
    InitHide(me : mutable)
	---C++: inline
    is static;
    
    MoreHide(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NextHide(me : mutable)
	---C++: inline
    is static;
    
    Hide(me : mutable; Coordinates : out Address    from Standard;
                       status      : out EdgeStatus from HLRAlgo;
		       S           : out Shape      from TopoDS;
                       reg1,regn   : out Boolean    from Standard;
                       outl,intl   : out Boolean    from Standard)
    is static;
    
    InitShow(me : mutable)
	---C++: inline
    is static;
    
    MoreShow(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    NextShow(me : mutable)
	---C++: inline
    is static;
    
    Show(me : mutable; Coordinates : out Address from Standard;
		       S           : out Shape   from TopoDS;
                       reg1,regn   : out Boolean from Standard;
                       outl,intl   : out Boolean from Standard)
    is static;
    
    OutLinedShape(me; S : Shape from TopoDS)
    returns Shape from TopoDS
	---Purpose: Make a shape  with  the internal outlines in  each
	--          face.
    is static;
    
    Debug(me) returns Boolean from Standard
	---C++: inline
    is static;
    
    Debug(me : mutable; B : Boolean from Standard)
	---C++: inline
    is static;
    
fields
    myProj       : Projector         from HLRAlgo;
    TMat         : Real              from Standard[3,3];
    TLoc         : Real              from Standard[3];
    TTMa         : Real              from Standard[3,3];
    TTLo         : Real              from Standard[3];
    TIMa         : Real              from Standard[3,3];
    TILo         : Real              from Standard[3];
    myShapes     : SequenceOfShape   from TopTools;
    myEMap       : IndexedMapOfShape from TopTools;
    myFMap       : IndexedMapOfShape from TopTools;
    myAlgo       : PolyAlgo          from HLRAlgo;
    myDebug      : Boolean           from Standard;
    myAngle      : Real              from Standard;
    myTolSta     : Real              from Standard;
    myTolEnd     : Real              from Standard;
    myTolAngular : Real              from Standard;
    myGSurf      : Surface           from Geom; 
    myBSurf      : Surface           from BRepAdaptor;
    myBCurv      : Curve             from BRepAdaptor;
    myPC         : Curve2d           from BRepAdaptor;

end PolyAlgo;
