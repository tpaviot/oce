-- Created on: 1995-10-10
-- Created by: GG
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class TransientManager from Visual3d inherits TShared

    ---Version:

    ---Purpose: This class allows to manage transient graphics
    --      above one View.
    --      A simple way to drawn something very quicly above
    --      a complex scene (Hilighting,Sketching,...)
    --      All transient graphics will be erased at the next
    --      View::BeginDraw().
    --      If RetainMode is active,
    --      All transient graphics will be kept at the
    --      next View::Update(),Redraw(). The transient graphics
    --      is stored by this object and graphic library, the 
    --      graphic managed itself exposure,resizing,...
    --      The method View::ClearDraw() is necessary to erase
    --      all transient graphics.
    --      If RetainMode is deactivate,
    --      All transient graphics will be erased at the
    --      next View::Update(),Redraw().
    --      Remember that nothing is stored by this object and
    --      graphic library,the application must managed itself
    --      exposure,resizing,...
    --      If double_buffering is activate,
    --      all graphics are drawn in the back buffer and flushed
    --      in the front buffer at the end of drawing but nothing
    --      is done for to separate transient from structured
    --      graphics,the only way to regenerate the structured
    --      view is to Redraw() the view.
    --      If double_buffering is deactivate,
    --      the back buffer is preserved and used for restoring 
    --      the front buffer at begin drawing time.I recommend
    --      to use the second way (without DB) if you want
    --      to preserve the graphics and the performances!
    
    
uses

    Array2OfReal             from TColStd,

    ExtendedString           from TCollection,

    PlaneAngle               from Quantity,

    Structure                from Graphic3d,
    AspectLine3d             from Graphic3d,
    AspectFillArea3d         from Graphic3d,
    AspectText3d             from Graphic3d,
    AspectMarker3d           from Graphic3d,
    TypeOfComposition        from Graphic3d,
    TextPath                 from Graphic3d,
    HorizontalTextAlignment  from Graphic3d,
    VerticalTextAlignment    from Graphic3d,

    View            from Visual3d

raises
    TransientDefinitionError from Visual3d,
    TransformError            from Graphic3d

is
    -------------------------
    -- Category: Constructors
    -------------------------

    Create returns mutable TransientManager from Visual3d;
    ---Purpose: Creates a TransientManager <aView>.
    ---Category: Constructors

    ------------------------
    -- Category: Destructors
    ------------------------

    Destroy (me : mutable);
    ---Level: Public
    ---Purpose: Suppress the TransientManager <me>.
    ---Category: Destructors
    ---C++: alias ~

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------

    BeginDraw (myclass;
           aView : View from Visual3d;
           DoubleBuffer: Boolean = Standard_False;
           RetainMode: Boolean = Standard_False)
    returns Integer from Standard
    ---Level: Public
    ---Purpose: Begins any graphics in the view <aView>
    --      Redraw any structured graphics in the back buffer before
    --      if <DoubleBuffer> is TRUE.
    --          Restore the front buffer from the back before
    --      if <DoubleBuffer> is FALSE.
    --      if <RetainMode> is TRUE.
    --          the graphic managed itself exposure,resizing ...
    --      if <RetainMode> is FALSE.
    --          the application must managed itself exposure,resizing ...
    --  
    --  Warning: Returns TRUE if transient drawing is enabled in
    --     the associated view.
    --          Returns FALSE ,if nothing works because something
    --     is wrong for the transient principle :
    --     Immediat mode is not implemented depending of the
    --     graphic library used.
    --         MBX,PIXMAP double buffering don't works depending of
    --         the graphic board and the visual of the window supporting 
    --         the view.
    --  Warning: No default attributes
    -- Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is already opened.
    -- or   the associated view is not mapped on a window.
    raises TransientDefinitionError from Visual3d;

    EndDraw (myclass;
         Synchronize: Boolean = Standard_False)
    ---Level: Public
    ---Purpose: Flush all graphics to the front buffer.
    --  Synchronize graphics to the screen if <Synchronize> is
    --  TRUE (make becarefull to the performances!).
        --  Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is not opened.
    raises TransientDefinitionError from Visual3d;

    ClearDraw (myclass; aView : View from Visual3d; 
                            aFlush : Boolean from Standard = Standard_True)
    ---Level: Public
    ---Purpose: Clear all transient graphics in the view <aView>
    ---         updates a scene if <aFlush> = true
        --  Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is already opened.
    -- or   the associated view is not mapped on a window.
    raises TransientDefinitionError from Visual3d;

    ---------------------------------------------------
    -- Category: Methods to modify the class definition
    ---------------------------------------------------

    BeginAddDraw (myclass;
           aView : View from Visual3d)
    returns Integer from Standard
    ---Level: Public
    ---Purpose: Begins any add graphics in the view <aView>
    --          the application must managed itself exposure,resizing ...
    --  
    --  Warning: Returns TRUE if transient drawing is enabled in
    --     the associated view.
    --          Returns FALSE ,if nothing works because something
    --     is wrong for the transient principle :
    --     Immediat mode is not implemented depending of the
    --     graphic library used.
    --         MBX,PIXMAP double buffering don't works depending of
    --         the graphic board and the visual of the window supporting 
    --         the view.
    --  Warning: No default attributes
        -- Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is already opened.
    -- or   the associated view is not mapped on a window.
    raises TransientDefinitionError from Visual3d;

    EndAddDraw (myclass)
    ---Purpose: Flush all add graphics to the front buffer.
    -- Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is not opened.
    raises TransientDefinitionError from Visual3d;

    ---------------------------------------
    -- Category: Graphic definition methods
    ---------------------------------------

    DrawStructure (myclass;
                AStructure   : Structure from Graphic3d)
        ---Purpose: Drawn the structure <AStructure>.
    -- Raises TransientDefinitionError from Visual3d;
    -- if   Drawing is not opened.
    raises TransientDefinitionError from Visual3d;

end TransientManager from Visual3d;
