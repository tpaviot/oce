-- Created on: 1997-04-17
-- Created by: Christophe MARION
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceData from HLRBRep

uses
    Boolean     from Standard,
    ShortReal   from Standard,
    Orientation from TopAbs,
    WiresBlock  from HLRAlgo,
    Surface     from HLRBRep,
    Face        from TopoDS

is
    Create returns FaceData from HLRBRep;

    Set(me : in out; FG  : Face        from TopoDS;
	             Or  : Orientation from TopAbs;
                     Cl  : Boolean     from Standard;
                     NW  : Integer     from Standard)
    	---Purpose: <Or> is the orientation of the face.  <Cl> is true
    	--          if the face  belongs to a  closed  volume. <NW> is
    	--          the number of wires ( or block  of  edges ) of the
    	--          face.
    is static;
    
    SetWire(me : in out; WI : Integer from Standard;
    	    	    	 NE : Integer from Standard)
    	---Purpose: Set <NE> the number  of  edges of the wire  number
    	--          <WI>.
    is static;
    
    SetWEdge(me : in out; WI,EWI,EI           : Integer     from Standard;
			  Or                  : Orientation from TopAbs;
                          OutL,Inte,Dble,IsoL : Boolean     from Standard)
    	---Purpose: Set the edge number <EWI> of the  wire <WI>.
    is static;
    
    Selected(me) returns Boolean from Standard
    	---C++: inline
    is static;
    
    Selected(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;
    
    Back(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Back(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Side(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Side(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Closed(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Closed(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Hiding(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Hiding(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Simple(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Simple(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Cut(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Cut(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    WithOutL(me) returns Boolean from Standard
    	---C++: inline
    is static;

    WithOutL(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Plane(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Plane(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Cylinder(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Cylinder(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Cone(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Cone(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Sphere(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Sphere(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Torus(me) returns Boolean from Standard
    	---C++: inline
    is static;

    Torus(me : in out; B : Boolean from Standard)
    	---C++: inline
    is static;

    Size(me) returns Real from Standard
    	---C++: inline
    is static;

    Size(me : in out; S : Real from Standard)
    	---C++: inline
    is static;

    Orientation(me) returns Orientation from TopAbs
        ---C++: inline
    is static;

    Orientation(me : in out; O : Orientation from TopAbs)
        ---C++: inline
    is static;

    Wires(me : in out) returns WiresBlock from HLRAlgo
        ---C++: inline
        ---C++: return &
    is static;

    Geometry(me : in out) returns Surface from HLRBRep
        ---C++: inline
        ---C++: return &
    is static;

    Tolerance(me) returns ShortReal from Standard
        ---C++: inline
    is static;

fields
    myFlags       : Integer    from Standard;
    myWires       : WiresBlock from HLRAlgo;
    myGeometry    : Surface    from HLRBRep;
    mySize        : Real       from Standard;
    myTolerance   : ShortReal  from Standard;

end FaceData;
