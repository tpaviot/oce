-- Created on: 1992-09-11
-- Created by: Stephan GARNAUD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EnvironmentIterator from OSD   

 ---Purpose: This allows consultation of every environment variable.
 --          There is no specific order of results.

uses Environment, Error, AsciiString from TCollection
raises OSDError

is
 Create returns EnvironmentIterator;
    ---Purpose: Instantiates Object as Iterator;
    ---Level: Public

 Destroy ( me : out );
	---C++: alias ~
	-- Only implemented on Windows NT system

 More (me : in out) returns Boolean  is static;
    ---Purpose: Returns TRUE if there are other environment variables.
    ---Level: Public

 Next (me : in out)  is static;
    ---Purpose: Sets the iterator to the next item.
    --          Returns the item value corresponding to the current
    --          position of the iterator.
    ---Level: Public

 Values (me : in out) returns Environment is static;
    ---Purpose: Returns the next environment variable found.
    ---Level: Public

 Failed (me) returns Boolean is static;
   ---Purpose: Returns TRUE if an error occurs
    ---Level: Public

 Reset (me : in out) is static;
   ---Purpose: Resets error counter to zero
    ---Level: Public
      
 Perror (me : in out)
   ---Purpose: Raises OSD_Error
    ---Level: Public
   raises OSDError is static ;

 Error (me) returns Integer is static ;
   ---Purpose: Returns error number if 'Failed' is TRUE.
    ---Level: Public

 fields
      myEnv        : Address;         -- Windows NT specific
      myCount      : CString;         -- Count in list of variables
      myError      : Error;
end EnvironmentIterator from OSD;

