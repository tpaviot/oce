-- Created on: 1992-11-17
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DispGlobal  from IFSelect  inherits Dispatch

    ---Purpose : A DispGlobal gathers all the input Entities into only one
    --           global Packet

uses AsciiString from TCollection, Graph, SubPartsIterator

is

    Create returns mutable DispGlobal;
    ---Purpose : Creates a DispGlobal

    Label (me) returns AsciiString from TCollection;
    ---Purpose : Returns as Label, "One File for all Input"

    	--  --    Evaluation    --  --

    LimitedMax (me; nbent : Integer; max : out Integer) returns Boolean
    	is redefined;
    ---Purpose : Returns True : maximum equates 1

    PacketsCount (me; G : Graph; count : out Integer) returns Integer
    	is redefined;
    ---Purpose : Returns True (count of packets is well known) and count is 1

    Packets (me; G : Graph; packs : in out SubPartsIterator);
    ---Purpose : Computes the list of produced Packets. It is made of only ONE
    --           Packet, which gets the RootResult from the Final Selection.
    --           Remark : the inherited exception raising is never activated.

end DispGlobal;
